module Frame_Buffer(output reg s,input a,input r0,input r1,input r2,input r3,input r4,input r5,input r6,input r7,input r8,input r9,input r10,input r11,input r12,input r13,input r14,input r15);
	
	reg [8:0] mem [80][30];
	
	
endmodule
