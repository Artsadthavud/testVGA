module Frame_Buffer(output reg s,input a);
	reg [10:0] mem [420];
endmodule
