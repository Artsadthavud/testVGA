module Frame_Buffer(output reg s,input a);
	
endmodule
